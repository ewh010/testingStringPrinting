//Group Name: 
//March 1, 2018
//This file will contain pipelining instructions: Fetch Decode Execute Mem Writeback


/********************** FETCH MODULE ***************************/
module Fetch(input [31:0] currPC, input [31:0] stall, output [31:0] PCF)

endmodule

/********************** DECODE MODULE ***************************/
module Decode(input [31:0] instr, output [31:0] instrD)

endmodule


/********************** EXECUTE MODULE ***************************/
module Execute()

endmodule

/********************** MEMORY MODULE ***************************/
module Mem()

endmodule

/********************** WRITEBACK MODULE ***************************/
module Writeback()
endmodule