//Group Name: 
//March 1, 2018
//This file will contain pipelining instructions: Fetch Decode Execute Mem Writeback


/********************** FETCH MODULE ***************************/
module Fetch(input [31:0] currPC, input [/*not sure how large*/] stallF, output [31:0]/*this is an assumption*/ PCF)

endmodule

/********************** DECODE MODULE ***************************/
module Decode(input [31:0] instr, input [/*not sure how large*/ ] stallD, output [31:0]/*this is an assumption*/ instrD)

endmodule


/********************** EXECUTE MODULE ***************************/
module Execute()

endmodule

/********************** MEMORY MODULE ***************************/
module Mem()

endmodule

/********************** WRITEBACK MODULE ***************************/
module Writeback()
endmodule